`include "constants.sv"
`include "registerfile.sv"
`include "alu.sv"
`include "controlpath.sv"