`include "datapath.sv"